library verilog;
use verilog.vl_types.all;
entity MSXPi_vlg_vec_tst is
end MSXPi_vlg_vec_tst;
