
rm  hardware/CPLD\ Project/*.done
rm  hardware/CPLD\ Project/*.jdi
rm  hardware/CPLD\ Project/db/*.cdb
rm  hardware/CPLD\ Project/db/*.hdb
rm  hardware/CPLD\ Project/db/*.qmsg
rm  hardware/CPLD\ Project/db/*.rdb
rm  hardware/CPLD\ Project/db/*.ddb
rm  hardware/CPLD\ Project/db/*.tdb
rm  hardware/CPLD\ Project/db/*.hif