library ieee;
use ieee.std_logic_1164.all;

package MSXPi_package is

        constant CTRLPORT1: STD_LOGIC_VECTOR(7 downto 0) := x"56";
        constant DATAPORT1: STD_LOGIC_VECTOR(7 downto 0) := x"5A";

end MSXPi_package;
